--Instruction decoder by Jakob & Yousef

-- library declaration
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;            -- basic IEEE library
use IEEE.NUMERIC_STD.ALL;               -- IEEE library for the unsigned type
                                        -- and various arithmetic operations

-- entity
entity inst_set is
	 
end inst_set;

-- architecture
architecture Behavioral of inst_set is



end Behavioral;

