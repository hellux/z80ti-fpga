library ieee;
use ieee.std_logic_1164.all;
use work.cmp_comm.all;
use work.z80_comm.all;
use work.ti_comm.all;

entity comp is port(
    clk : in std_logic;
-- dbg input
    btns : in std_logic_vector(4 downto 0);
    sw : in std_logic_vector(7 downto 0);
-- keyboard
    ps2_kbd_clk : in std_logic;
    ps2_kbd_data : in std_logic;
-- vga monitor
    vga_red : out std_logic_vector(2 downto 0);
    vga_green : out std_logic_vector(2 downto 0);
    vga_blue : out std_logic_vector(2 downto 1);
    hsync, vsync : out std_logic;
-- memory
    maddr : out std_logic_vector(25 downto 0);
    mdata : inout std_logic_vector(15 downto 0);
    mclk, madv_c, mcre, mce_c, moe_c, mwe_c : out std_logic;
    mlb_c, mub_c : out std_logic;
-- 7 segment, led
    seg, led : out std_logic_vector(7 downto 0);
    an : out std_logic_vector(3 downto 0));
end comp;

architecture arch of comp is
    component z80 port(
        clk, ce : in std_logic;
        cbi : in ctrlbus_in;
        cbo : out ctrlbus_out;
        addr : out std_logic_vector(15 downto 0);
        data_in : in std_logic_vector(7 downto 0);
        data_out : out std_logic_vector(7 downto 0);
        dbg : out dbg_z80_t);
    end component;

    component ti port(
        clk, rst : in std_logic;
        int : out std_logic;
        cbo : in ctrlbus_out;
        addr_log : in std_logic_vector(15 downto 0);
        data_in : in std_logic_vector(7 downto 0);
        data_out : out std_logic_vector(7 downto 0);
        keys_down : in keys_down_t;
        on_key_down : in std_logic;
        x_vga : in std_logic_vector(6 downto 0);
        y_vga : in std_logic_vector(5 downto 0);
        data_vga : out std_logic;
        rd, wr : out std_logic;
        addr_phy : out std_logic_vector(19 downto 0));
    end component;

    component mem_if port(
        clk, rst : in std_logic;
        rd, wr : in std_logic;
        addr_phy : in std_logic_vector(19 downto 0);
        data_in : in std_logic_vector(7 downto 0);
        data_out : out std_logic_vector(7 downto 0);
    -- external
        maddr : out std_logic_vector(25 downto 0);
        mdata : inout std_logic_vector(15 downto 0);
        mclk, madv_c, mcre, mce_c, moe_c, mwe_c : out std_logic;
        mlb_c, mub_c : out std_logic);
    end component;

    component vga_motor port(
         clk : in std_logic;
         data : in std_logic;
         rst : in std_logic;
         x : out std_logic_vector(6 downto 0);
         y : out std_logic_vector(5 downto 0);
         vgaRed	: out std_logic_vector(2 downto 0);
         vgaGreen : out std_logic_vector(2 downto 0);
         vgaBlue : out std_logic_vector(2 downto 1);
         Hsync : out std_logic;
         Vsync : out std_logic);
    end component;

    component kbd_enc port (
        clk, rst : in std_logic;
        PS2KeyboardCLK : in std_logic;
        PS2KeyboardData	: in std_logic;
        keys_down : out keys_down_t;
        on_key_down : out std_logic;
        scancode_out : out std_logic_vector(7 downto 0);
        keycode_out : out std_logic_vector(7 downto 0));
    end component;

    component memory port(
        clk, rst : in std_logic;
        cbo : in ctrlbus_out;
        addr : in std_logic_vector(15 downto 0);
        data_in : in std_logic_vector(7 downto 0);
        data_out : out std_logic_vector(7 downto 0));
    end component;

    component monitor port(
        clk : in std_logic;
        sw : in std_logic_vector(5 downto 0);
        dbg : in dbg_cmp_t;
        seg, led : out std_logic_vector(7 downto 0);
        an : out std_logic_vector(3 downto 0));
    end component;

    constant DIV_6MHZ : integer := 17;
    constant DIV_TI : integer := 2;
    constant DIV_10HZ : integer := 10*10**6;
    constant DIV_100HZ : integer := 10**6;

    signal clk_cpu, clk_6mhz, clk_ti, clk_10hz, clk_100hz: std_logic;
    signal clk_6mhz_div : integer range 0 to DIV_6MHZ-1;
    signal clk_ti_div : integer range 0 to DIV_TI-1;
    signal clk_10hz_div : integer range 0 to DIV_10HZ-1;
    signal clk_100hz_div : integer range 0 to DIV_100HZ-1;

    signal cbo : ctrlbus_out;
    signal addr : std_logic_vector(15 downto 0);
    signal cbi : ctrlbus_in;
    signal int : std_logic;
    signal data, data_z80, data_mem, data_ti : std_logic_vector(7 downto 0);

    signal rst : std_logic;

    signal btns_sync, btns_q, btns_op : std_logic_vector(4 downto 0);

    signal dbg : dbg_cmp_t;

    -- ti <-> kbd
    signal keys_down : keys_down_t;
    signal on_key_down : std_logic := '0';
    -- ti <-> vga
    signal data_vga : std_logic;
    signal x_vga : std_logic_vector(6 downto 0);
    signal y_vga : std_logic_vector(5 downto 0);
    -- ti <-> mem controller
    signal mem_rd, mem_wr : std_logic;
    signal addr_phy : std_logic_vector(19 downto 0);
begin
    -- input sync
    op_btns : process(clk) begin
        if rising_edge(clk) then
            btns_sync <= btns;
            btns_q <= btns_sync;
        end if;
    end process;
    btns_op <= btns_sync and not btns_q;

    -- clock sync
    process(clk) begin
        if rising_edge(clk) then
            if clk_6mhz_div = DIV_6MHZ-1 then
                clk_6mhz_div <= 0;
            else
                clk_6mhz_div <= clk_6mhz_div + 1;
            end if;
            if clk_ti_div = DIV_TI-1 then
                clk_ti_div <= 0;
            else
                clk_ti_div <= clk_ti_div + 1;
            end if;
            if clk_10hz_div = DIV_10HZ-1 then
                clk_10hz_div <= 0;
            else
                clk_10hz_div <= clk_10hz_div + 1;
            end if;
            if clk_100hz_div = DIV_100HZ-1 then
                clk_100hz_div <= 0;
            else
                clk_100hz_div <= clk_100hz_div + 1;
            end if;
            if rst = '1' then
                clk_6mhz_div <= 0;
                clk_ti_div <= 0;
                clk_10hz_div <= 0;
                clk_100hz_div <= 0;
            end if;
        end if;
    end process;
    clk_6mhz  <= '1' when clk_6mhz_div  = 0 else '0';
    clk_ti    <= '1' when clk_ti_div    = 0 else '0';
    clk_100hz <= '1' when clk_100hz_div = 0 else '0';
    clk_10hz  <= '1' when clk_10hz_div  = 0 else '0';
    with sw(7 downto 6) select
        clk_cpu <= clk_100hz  when "01",
                   clk_10hz   when "10",
                   btns_op(0) when "11",
                   clk_6mhz   when others;

    -- buses
    rst <= btns(1);
    cbi.wt <= '0';
    cbi.int <= int;
    cbi.reset <= rst;
    -- OR data bus instead of tristate
    data <= data_z80 or data_mem or data_ti;

    -- cpu / asic
    cpu : z80 port map(clk, clk_cpu, cbi, cbo, addr, data, data_z80, dbg.z80);
    ti_comp : ti port map(clk_ti, rst,
                          int, cbo, addr, data, data_ti,
                          keys_down, on_key_down,
                          x_vga, y_vga, data_vga,
                          mem_rd, mem_wr, addr_phy);

    -- external controllers
    vga : vga_motor port map(clk, data_vga, rst, x_vga, y_vga,
                             vga_red, vga_green, vga_blue, hsync, vsync);
    mif : mem_if port map(clk, rst, mem_rd, mem_wr, addr_phy, data, data_mem,
                          maddr, mdata, mclk, madv_c, mcre, mce_c, moe_c,
                          mwe_c, mlb_c, mub_c);
    kbd : kbd_enc port map(clk, rst, ps2_kbd_clk, ps2_kbd_data,
                           keys_down, on_key_down, dbg.scancode, dbg.keycode);

    -- debug
    dbg.mem_rd <= mem_rd;
    dbg.mem_wr <= mem_wr;
    dbg.on_key_down <= on_key_down;
    dbg.data <= data;
    dbg.data_mem <= data_mem;
    dbg.addr_log <= addr;
    dbg.data_mem <= data_mem;
    dbg.addr_phy <= addr_phy;
    dbg.cbi <= cbi;
    dbg.cbo <= cbo;

    mon : monitor port map(clk, sw(5 downto 0), dbg, seg, led, an);
end arch;
